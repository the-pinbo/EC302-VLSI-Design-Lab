magic
tech scmos
timestamp 1667136153
<< nwell >>
rect -29 -18 60 42
<< polysilicon >>
rect -1 15 3 17
rect 12 15 16 17
rect 27 15 31 17
rect -1 -49 3 0
rect 12 -49 16 0
rect 27 -49 31 0
rect -1 -58 3 -56
rect 12 -58 16 -56
rect 27 -58 31 -56
<< ndiffusion >>
rect -9 -53 -7 -49
rect -3 -53 -1 -49
rect -9 -56 -1 -53
rect 3 -56 12 -49
rect 16 -52 27 -49
rect 16 -56 20 -52
rect 24 -56 27 -52
rect 31 -53 37 -49
rect 31 -56 41 -53
<< pdiffusion >>
rect -9 4 -1 15
rect -9 0 -7 4
rect -3 0 -1 4
rect 3 11 5 15
rect 9 11 12 15
rect 3 0 12 11
rect 16 4 27 15
rect 16 0 20 4
rect 24 0 27 4
rect 31 4 41 15
rect 31 0 37 4
<< metal1 >>
rect -5 33 -3 37
rect 1 33 5 37
rect 9 33 33 37
rect 37 33 40 37
rect 5 15 9 33
rect -7 -5 -3 0
rect 20 -5 24 0
rect -7 -9 24 -5
rect 37 -33 41 0
rect -7 -37 41 -33
rect -7 -49 -3 -37
rect 37 -49 41 -37
rect 20 -73 24 -56
rect -11 -74 45 -73
rect -11 -78 -9 -74
rect -5 -78 20 -74
rect 24 -78 37 -74
rect 41 -78 45 -74
<< ntransistor >>
rect -1 -56 3 -49
rect 12 -56 16 -49
rect 27 -56 31 -49
<< ptransistor >>
rect -1 0 3 15
rect 12 0 16 15
rect 27 0 31 15
<< polycontact >>
rect -5 -27 -1 -23
rect 8 -27 12 -23
rect 23 -27 27 -23
<< ndcontact >>
rect -7 -53 -3 -49
rect 20 -56 24 -52
rect 37 -53 41 -49
<< pdcontact >>
rect -7 0 -3 4
rect 5 11 9 15
rect 20 0 24 4
rect 37 0 41 4
<< psubstratepcontact >>
rect -9 -78 -5 -74
rect 20 -78 24 -74
rect 37 -78 41 -74
<< nsubstratencontact >>
rect -3 33 1 37
rect 5 33 9 37
rect 33 33 37 37
<< labels >>
rlabel metal1 15 34 15 34 1 vdd
rlabel polycontact -3 -25 -3 -25 1 a
rlabel polycontact 10 -25 10 -25 1 b
rlabel polycontact 25 -25 25 -25 1 c
rlabel metal1 14 -76 14 -76 1 vss
rlabel metal1 39 -26 39 -26 1 vout
<< end >>
