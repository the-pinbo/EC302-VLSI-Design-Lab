magic
tech scmos
timestamp 1667131608
<< nwell >>
rect -14 9 12 43
<< polysilicon >>
rect -6 32 -4 34
rect 2 32 4 34
rect -6 6 -4 22
rect 2 6 4 22
rect -10 2 -4 6
rect -2 2 4 6
rect -6 -2 -4 2
rect 2 -2 4 2
rect -6 -9 -4 -7
rect 2 -9 4 -7
<< ndiffusion >>
rect -11 -3 -6 -2
rect -7 -7 -6 -3
rect -4 -7 2 -2
rect 4 -6 5 -2
rect 4 -7 9 -6
<< pdiffusion >>
rect -11 29 -6 32
rect -7 25 -6 29
rect -11 22 -6 25
rect -4 29 2 32
rect -4 25 -3 29
rect 1 25 2 29
rect -4 22 2 25
rect 4 29 9 32
rect 4 25 5 29
rect 4 22 9 25
<< metal1 >>
rect -6 36 4 41
rect -3 29 1 36
rect -11 14 -7 25
rect 5 14 9 25
rect -11 10 9 14
rect 5 -2 9 10
rect -11 -13 -7 -7
rect -6 -18 4 -13
<< ntransistor >>
rect -6 -7 -4 -2
rect 2 -7 4 -2
<< ptransistor >>
rect -6 22 -4 32
rect 2 22 4 32
<< ndcontact >>
rect -11 -7 -7 -3
rect 5 -6 9 -2
<< pdcontact >>
rect -11 25 -7 29
rect -3 25 1 29
rect 5 25 9 29
<< psubstratepcontact >>
rect -11 -18 -6 -13
rect 4 -18 9 -13
<< nsubstratencontact >>
rect -11 36 -6 41
rect 4 36 9 41
<< labels >>
rlabel metal1 -1 38 -1 38 1 vdd
rlabel polysilicon -8 4 -8 4 7 a
rlabel polysilicon 0 4 0 4 7 b
rlabel metal1 7 4 7 4 3 out
rlabel metal1 -1 -16 -1 -16 5 vss
<< end >>
