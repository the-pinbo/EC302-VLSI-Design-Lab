magic
tech scmos
timestamp 1667378637
<< nwell >>
rect -5 -4 27 25
<< polysilicon >>
rect 3 14 7 16
rect 15 14 19 16
rect 3 -13 7 -1
rect 15 -13 19 -1
rect 3 -30 7 -28
rect 15 -30 19 -28
<< ndiffusion >>
rect -5 -19 3 -13
rect -5 -23 -3 -19
rect 1 -23 3 -19
rect -5 -28 3 -23
rect 7 -28 15 -13
rect 19 -17 21 -13
rect 25 -17 27 -13
rect 19 -28 27 -17
<< pdiffusion >>
rect -5 4 3 14
rect -5 0 -3 4
rect 1 0 3 4
rect -5 -1 3 0
rect 7 12 15 14
rect 7 8 9 12
rect 13 8 15 12
rect 7 -1 15 8
rect 19 4 27 14
rect 19 0 21 4
rect 25 0 27 4
rect 19 -1 27 0
<< metal1 >>
rect -5 32 27 33
rect -5 28 9 32
rect 13 28 27 32
rect -5 25 27 28
rect 9 12 13 25
rect 1 0 21 4
rect 21 -5 25 0
rect 21 -9 29 -5
rect 21 -13 25 -9
rect -3 -32 1 -23
rect -5 -34 27 -32
rect -5 -38 9 -34
rect 13 -38 27 -34
rect -5 -40 27 -38
<< ntransistor >>
rect 3 -28 7 -13
rect 15 -28 19 -13
<< ptransistor >>
rect 3 -1 7 14
rect 15 -1 19 14
<< polycontact >>
rect -1 -11 3 -7
rect 11 -11 15 -7
<< ndcontact >>
rect -3 -23 1 -19
rect 21 -17 25 -13
<< pdcontact >>
rect -3 0 1 4
rect 9 8 13 12
rect 21 0 25 4
<< psubstratepcontact >>
rect 9 -38 13 -34
<< nsubstratencontact >>
rect 9 28 13 32
<< labels >>
rlabel metal1 -5 33 27 33 1 vdd
rlabel polycontact -1 -11 -1 -7 7 v_a
rlabel metal1 -5 -40 27 -40 1 vss
rlabel polycontact 11 -11 11 -7 1 v_b
rlabel metal1 29 -9 29 -5 7 vout
<< end >>
