magic
tech scmos
timestamp 1667379706
<< polysilicon >>
rect -22 55 -18 57
rect -10 55 -6 57
rect 19 46 23 49
rect -22 27 -18 39
rect -10 27 -6 39
rect 19 34 23 38
rect 9 30 23 34
rect 19 26 23 30
rect -22 21 -18 23
rect -10 21 -6 23
rect 19 19 23 22
<< ndiffusion >>
rect -24 23 -22 27
rect -18 23 -16 27
rect -12 23 -10 27
rect -6 23 -4 27
rect 15 22 19 26
rect 23 22 27 26
<< pdiffusion >>
rect -24 51 -22 55
rect -28 39 -22 51
rect -18 39 -10 55
rect -6 47 0 55
rect -6 42 -5 47
rect -6 39 0 42
rect 15 42 19 46
rect 11 38 19 42
rect 23 42 31 46
rect 23 38 27 42
<< metal1 >>
rect -28 73 32 74
rect -28 69 -16 73
rect -12 69 32 73
rect -28 66 32 69
rect -28 55 -24 66
rect -16 59 8 62
rect -16 47 -12 59
rect -16 42 -5 47
rect -16 27 -12 42
rect 5 34 8 59
rect 11 46 15 66
rect 27 26 31 38
rect -28 8 -24 23
rect -4 8 0 23
rect 11 8 15 22
rect -28 6 32 8
rect -28 2 -16 6
rect -12 2 32 6
rect -28 0 32 2
<< ntransistor >>
rect -22 23 -18 27
rect -10 23 -6 27
rect 19 22 23 26
<< ptransistor >>
rect -22 39 -18 55
rect -10 39 -6 55
rect 19 38 23 46
<< polycontact >>
rect -26 30 -22 34
rect -6 34 -2 38
rect 5 30 9 34
<< ndcontact >>
rect -28 23 -24 27
rect -16 23 -12 27
rect -4 23 0 27
rect 11 22 15 26
rect 27 22 31 26
<< pdcontact >>
rect -28 51 -24 55
rect -5 42 0 47
rect 11 42 15 46
rect 27 38 31 42
<< psubstratepcontact >>
rect -16 2 -12 6
<< nsubstratencontact >>
rect -16 69 -12 73
<< labels >>
rlabel metal1 -28 74 0 74 1 vdd
rlabel polycontact -26 30 -26 34 3 v_a
rlabel metal1 -28 0 0 0 5 vss
rlabel polycontact -2 34 -2 38 7 v_b
rlabel metal1 29 32 29 32 3 vout
<< end >>
